module controller(

); 

endmodule