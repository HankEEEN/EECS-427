`timescale 1ns/1ps

`ifndef CLK_PERIOD
 `define CLK_PERIOD 20
`endif

module pc_nop_tb;

parameter   ADDR_WIDTH = 16;
parameter   DISP_WIDTH = 8;





endmodule